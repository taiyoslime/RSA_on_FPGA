
`define mbit 63;
`define mbit_h 31;
